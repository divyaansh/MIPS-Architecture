library verilog;
use verilog.vl_types.all;
entity tb_8bit2to1mux is
end tb_8bit2to1mux;
